// Copyright 2021 Datum Technology Corporation
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
// Licensed under the Solderpad Hardware License v 2.1 (the "License"); you may not use this file except in compliance
// with the License, or, at your option, the Apache License version 2.0.  You may obtain a copy of the License at
//                                        https://solderpad.org/licenses/SHL-2.1/
// Unless required by applicable law or agreed to in writing, any work distributed under the License is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_AXIS_IF_CHKR_SV__
`define __UVMA_AXIS_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_axis_if.
 */
module uvma_axis_if_chkr(
   uvma_axis_if  axis_if
);
   
   // TODO Add assertions to uvma_axis_if_chkr
   
endmodule : uvma_axis_if_chkr


`endif // __UVMA_AXIS_IF_CHKR_SV__
