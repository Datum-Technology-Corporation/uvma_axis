// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_AXIS_ST_MACROS_SV__
`define __UVMT_AXIS_ST_MACROS_SV__


`ifndef UVMT_AXIS_ST_CLI_ARG_NUM_TRANSFERS
   `define UVMT_AXIS_ST_CLI_ARG_NUM_TRANSFERS "NTRN"
`endif
`ifndef UVMT_AXIS_ST_CLI_ARG_MIN_TRANSFER_SIZE
   `define UVMT_AXIS_ST_CLI_ARG_MIN_TRANSFER_SIZE "MINSZ"
`endif
`ifndef UVMT_AXIS_ST_CLI_ARG_MAX_TRANSFER_SIZE
   `define UVMT_AXIS_ST_CLI_ARG_MAX_TRANSFER_SIZE "MAXSZ"
`endif
`ifndef UVMT_AXIS_ST_CLI_ARG_MIN_GAP
   `define UVMT_AXIS_ST_CLI_ARG_MIN_GAP "MINGAP"
`endif
`ifndef UVMT_AXIS_ST_CLI_ARG_MAX_GAP
   `define UVMT_AXIS_ST_CLI_ARG_MAX_GAP "MAXGAP"
`endif
`ifndef UVMT_AXIS_ST_CLI_ARG_MSTR_TON
   `define UVMT_AXIS_ST_CLI_ARG_MSTR_TON "MSTRON"
`endif
`ifndef UVMT_AXIS_ST_CLI_ARG_SLV_TON
   `define UVMT_AXIS_ST_CLI_ARG_SLV_TON "SLVON"
`endif


`endif // __UVMT_AXIS_ST_MACROS_SV__
