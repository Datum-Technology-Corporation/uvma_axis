// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_AXIS_ST_CHKR_SV__
`define __UVME_AXIS_ST_CHKR_SV__


/**
 * TODO Describe uvme_axis_st_chkr
 */
module uvme_axis_st_chkr (
      uvma_axis_if  mstr_if,
      uvma_axis_if  slv_if
);
   
   // TODO Add assertions to uvme_axis_st_chkr
   
endmodule : uvme_axis_st_chkr


`endif // __UVME_AXIS_ST_CHKR_SV__
