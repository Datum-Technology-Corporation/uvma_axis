// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_AXIS_ST_BASE_TEST_WORKAROUNDS_SV__
`define __UVMT_AXIS_ST_BASE_TEST_WORKAROUNDS_SV__


// This file should be empty by the end of the project

constraint mstr_ton_cons {
   
}


`endif // __UVMT_AXIS_ST_BASE_TEST_WORKAROUNDS_SV__
