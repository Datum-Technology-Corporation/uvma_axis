// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_AXIS_ST_DUT_CHKR_SV__
`define __UVMT_AXIS_ST_DUT_CHKR_SV__


/**
 * Module encapsulating assertions for AMBA Advanced Extensible Interface Stream Agent Self-Testing DUT wrapper
 * (uvmt_axis_st_dut_wrap).
 */
module uvmt_axis_st_dut_chkr(
   uvma_axis_if  mstr_if,
   uvma_axis_if  slv_if
);
   
   // TODO Add assertions to uvmt_axis_st_dut_chkr
   
endmodule : uvmt_axis_st_dut_chkr


`endif // __UVMT_AXIS_ST_DUT_CHKR_SV__
