// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_AXIS_IF_CHKR_SV__
`define __UVMA_AXIS_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_axis_if.
 */
module uvma_axis_if_chkr (
   uvma_axis_if  axis_if
);
   
   // TODO Add assertions to uvma_axis_if_chkr
   
endmodule : uvma_axis_if_chkr


`endif // __UVMA_AXIS_IF_CHKR_SV__
